`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:15:49 11/18/2017 
// Design Name: 
// Module Name:    Simulation 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Simulation(input clk, output reg r
    );
reg[5131:0]E;
reg [683:0]A;
reg [341:0]B;
reg [41:0]T;
reg [41:0]D;
reg [5131:0]H;
integer w =5131;
integer cn=0;
integer leds=49;
integer q=0;
always@(posedge clk)
begin
if(q==654)
begin
	A=684'b1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_1000;
	B=342'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0;
	T=42'b1000_1000_1000_1000_1000_1000_1000_1000_1000_1000_10;
	D=42'b00000_00000_00000_00000_00000_00000_00000_00000_00000_00000_00;
	H=E;
	case(leds)
	112:E={A,B,T,D,T,D,T,D,D,D,T,D, T,D,T,D,T,D,T,D ,T,D,D,D, T,D,D,D, T,D,T,D,D,D ,T,D,D,D, T,D,D,D,T,D,D,D,T,D,D,D ,T,D,T,D,T,D,T,D,D,D ,T,D,T,D,T,D,T,D , T,D,D,D,T,D,D,D, T,D,D,D, T,D , T,D,D,D, T,D,D,D, T,D,D,D, T,D,D,D ,A[42:0]};

49:E={A,B,T,D,T,D,T,D,D,D,T,D, T,D,T,D,T,D,T,D ,T,D,D,D, T,D,D,D, T,D,T,D,D,D ,T,D,D,D, T,D,D,D,T,D,D,D,T,D,D,D ,T,D,D,D,T,D,T,D,T,D ,T,D,D,D,T,D,T,D,T,D , T,D,T,D,D,D, T,D,D,D, T,D,D,D , T,D,T,D,D,D, T,D,D,D, T,D,D,D ,A[42:0]};

50:E={A,B,T,D,T,D,T,D,D,D,T,D, T,D,T,D,T,D,T,D ,T,D,D,D, T,D,D,D, T,D,T,D,D,D ,T,D,D,D, T,D,D,D,T,D,D,D,T,D,D,D ,T,D,T,D,D,D,T,D,T,D ,T,D,D,D,T,D,T,D,T,D , T,D,D,D,T,D, T,D,D,D, T,D,D,D , T,D,T,D,D,D, T,D,D,D, T,D,D,D ,A[42:0]};

51:E={A,B,T,D,T,D,T,D,D,D,T,D, T,D,T,D,T,D,T,D ,T,D,D,D, T,D,D,D, T,D,T,D,D,D ,T,D,D,D, T,D,D,D,T,D,D,D,T,D,D,D ,T,D,D,D,T,D,D,D,T,D,T,D ,T,D,D,D,T,D,T,D,T,D , T,D,T,D, T,D,D,D, T,D,D,D , T,D,T,D,D,D, T,D,D,D, T,D,D,D ,A[42:0]};
endcase
	if(H!=E)
		cn=0;
	if(w>-1&&cn==0)
		begin
		r=E[w];
		w=w-1;
		end
	else
		begin
		r=0;
		w=5131;
		cn=1;
		end
q=0;
end
else q=q+1;
end
endmodule


